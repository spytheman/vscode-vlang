module main

fn main() {
	
}
